package WiredParam

// 后端允许的 Checkpoint/Branch Issue Queue 尺寸
typedef 4 BRANCH_SLOT


endpackage : WiredParam