// Wired 核心中，MTLB采用 FPGA 不友好的 CAM 电路实现;
// 因此尽量保持较低的规格，避免较大的组合逻辑导致频率过低。
// 按照设计，MTLB 中仅存储巨页（16M/8M），此 MTLB 仅需要支持 Linux 中存在的几种巨页配置即可
// 表项数维持在 4-16 项。
