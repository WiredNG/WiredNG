`ifndef _WIREDNG_BRANCH_HEADER_
`define _WIREDNG_BRANCH_HEADER_

`include "wiredng_params.svh"

typedef struct packed {
    logic[47:0]
} ftq_entry_t;

`endif