package WiredParam

// 后端允许的 Checkpoint/Branch Issue Queue 尺寸
typedef 4 BRANCH_SLOT

typedef 64 FP_PHYREG_NUM
typedef 64 INT_PHYREG_NUM

endpackage : WiredParam