// Wired 核心中，MTLB采用 FPGA 不友好的 CAM 电路实现;
// 因此尽量保持较低的规格，避免较大的组合逻辑导致频率过低。
