package Dividers;



endpackage : Dividers

