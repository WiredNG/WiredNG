// Wired 下一代核心模块：Load ROB