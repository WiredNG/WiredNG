package WiredDecode

import WiredTypes::*;
import WiredParam::*;

endpackage : WiredDecode