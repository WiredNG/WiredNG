// Wired 下一代核心，硬件页表遍历模块
// Wired 下一代核心采用 TLB 硬件重填实现，对于所有 TLB 缺失，进行硬件重填
// 注意：硬件 PTW 与 3A6000 中实现不一致，不支持 fast-path。PTW 对于内存是只读的。
// 仍需要软件维护 TLB 与内存页表的一致性，包括解决 TLB Shutdown 问题。

module wiredng_ptw (
    input wire clk,
    input wire rst_n,

    
);

endmodule