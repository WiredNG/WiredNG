// 下一代 Wired 核心， Commited store buffer
// Cache 内部模块，按写端口粒度组织
module wiredng_csb(
    input wire clk,
    input wire rst_n
);

endmodule