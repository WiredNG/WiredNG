// 前端取指队列
// 采用类似 ROB 的设计逻辑
// 由于取值部分存在乱序可能（靠后取指先写入）
// 因此取值队列内部也维护一个 id，由 id 完成读写。
// 有效性判断采用双寄存器堆 XOR 的方式实现